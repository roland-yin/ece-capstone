module controller #(
    parameter FRAC = 15
) (
    input  wire                 clk,
    input  wire                 rst_n,
    input  wire                 in_valid,       // from input_buffer
    input  wire signed [15:0]   e_in,
    input  wire signed [15:0]   x_in,
    input  wire signed [15:0]   a_in,
    input  wire signed [15:0]   u_in,           // step-size

    input  wire                 fir_done,       // FIR done signal
    input  wire signed [31:0]   fir_out,        // FIR output

    output reg  signed [15:0]   x_out,          // feed to FIR
    output reg  signed [15:0]   weight_adjust,  // (e - a) * u
    output reg  signed [31:0]   out_sample,     // core output from FIR
    output reg                  out_valid,      // core output ready
    output reg                  fir_go          // go signal for FIR
);

    reg signed [15:0] mult_a, mult_b;
    reg signed [31:0] mult_p;
    bw_mult bw_mult_weight_adjust (.a(mult_a), .b(mult_b), .p(mult_p));

    localparam S_IDLE = 2'd0, S_START = 2'd1, S_RUN = 2'd2, S_DONE = 2'd3;
    reg [1:0] state;

    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            state <= S_IDLE;
            x_out <= 32'sd0;
            weight_adjust <= 15'sd0;
            out_sample <= 32'sd0;
            out_valid <= 1'b0;
            fir_go <= 1'b0;
        end else begin
            out_valid <= 1'b0; // default
            fir_go <= 1'b0;    // default

            case (state)
                S_IDLE: begin
                    if (in_valid) begin
                        // compute weight adjustment
                        mult_a <= e_in - a_in;
                        mult_b <= u_in;
                        state <= S_START;
                    end
                end

                S_START: begin
                    weight_adjust <= mult_p;
                    x_out <= x_in;      // feed input to FIR
                    fir_go <= 1'b1;     // signal FIR to start
                    state <= S_RUN;
                end

                S_RUN: begin
                    // wait for FIR to finish
                    if (fir_done) begin
                        // capture FIR output
                        out_sample <= fir_out;
                        out_valid <= 1'b1;  // core output ready
                        state <= S_DONE;
                    end
                end

                S_DONE: begin
                    state <= S_IDLE; // ready for next input
                end
            endcase
        end
    end

endmodule
